** Profile: "SCHEMATIC1-time"  [ D:\scoala\an II\sem 2\computer aided design\project\project\project-pspicefiles\schematic1\time.sim ] 

** Creating circuit file "time.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\scoala\programe\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "D:\scoala\programe\Cadence\SPB_16.5\tools\pspice\library\nom.lib" 
.lib "D:\scoala\programe\Cadence\SPB_16.5\tools\pspice\library\nomd.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 SKIPBP 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
